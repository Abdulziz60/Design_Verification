
module top;

  // Instantiate the main testbench module
  router_tb tb();

endmodule
