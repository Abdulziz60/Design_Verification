interface dut_if ;
    
endinterface // 



