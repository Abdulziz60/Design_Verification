interface adder_if ;

    logic clk;
    logic [7:0] a, b , sum;
    logic Carry;

endinterface