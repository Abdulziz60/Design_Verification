module dut (dut_if aif);

endmodule