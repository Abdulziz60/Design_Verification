interface dut_if (input clk);
    logic [7:0] a;
    logic [7:0] b;
    logic [7:0] sum;
    logic carry;
endinterface // 



