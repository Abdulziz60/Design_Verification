module dut ( dut_if  dif);

endmodule