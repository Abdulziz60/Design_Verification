module TB;
initial begin
$display("Hello, SystemVerilog!");
end
endmodule
