
interface i2c_if (input logic clk);

    wire sda;
    wire scl;

endinterface