
`include "uvm_macros.svh"
import uvm_pkg::*;
import yapp_pkg::*;

module router_tb;

  initial begin
    run_test(); // runs base_test by default
  end

endmodule
