module top;
// import the UVM library
// include the UVM macros

// import the YAPP package

// generate 5 random packets and use the print method
// to display the results

// experiment with the copy, clone and compare UVM method
endmodule : top
