// Define your enumerated type(s) here

class yapp_packet extends uvm_sequence_item;

// Follow the lab instructions to create the packet.
// Place the packet declarations in the following order:

  // Define protocol data

  // Define control knobs

  // Enable automation of the packet's fields

  // Define packet constraints

  // Add methods for parity calculation and class construction

endclass: yapp_packet
